module lod_testbench;
  wire out;
  reg data_in;

  lod dut0(data
