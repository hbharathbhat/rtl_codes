module lod
